module resetar (A, S);

input  [3:0]A;
output  [3:0]S; 

assign S[0] = 0;
assign S[1] = 0;
assign S[2] = 0;
assign S[3] = 0;
 
endmodule